`include "uvm_macros.svh"
import uvm_pkg::*;
 
 
module tb;
  
  initial begin
    `uvm_info("TB_TOP","Hello_RTL",UVM_NONE);
  end
  
endmodule
